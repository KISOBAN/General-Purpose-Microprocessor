library verilog;
use verilog.vl_types.all;
entity FourtoSixteenDecoder_vlg_vec_tst is
end FourtoSixteenDecoder_vlg_vec_tst;
