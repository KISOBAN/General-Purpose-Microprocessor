LIBRARY IEEE;
USE ieee.std_logic_1164.all;
ENTITY FLIPFLOP IS
	PORT (
			 D : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			 CLK : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			 Q   : OUT STD_LOGIC VECTOR (1 DOWNTO 0));
END FLIPFLOP;
ARCHITECTURE BEHAVIOUR OF FLIPFLOP IS
	 signal Qreg : STD_LOGIC_VECTOR (1 DOWNTO 0);
BEGIN
PROCESS (D, CLK, Qreg)
BEGIN
			IF (CLK = '0') THEN
				Qreg <= Qreg;
			ELSIF (CLK'EVENT AND CLK = '1') THEN
				Qreg <= D;
			END IF;
END PROCESS;
Q <= Qreg;
END BEHAVIOUR;
				
			