library verilog;
use verilog.vl_types.all;
entity Lab6block_vlg_vec_tst is
end Lab6block_vlg_vec_tst;
